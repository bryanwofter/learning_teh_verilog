module draw_driver_core#(
    parameter SIZE = 1
) (
    input wire clk,
    input wire enable
);

endmodule
